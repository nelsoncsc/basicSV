interface four_bits_output_if();
  logic [3:0] c;
  modport port(output c);
endinterface: four_bits_output_if
