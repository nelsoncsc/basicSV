interface one_bit_input_if(input logic a, b);
  logic a, b;
  modport port(input a, b);
endinterface: one_bit_input_if
