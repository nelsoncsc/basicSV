interface four_bits_input_if(input logic[3:0] a, b);
  logic [3:0] a, b;
  modport port(input a, b);
endinterface: four_bits_input_if
