interface one_bit_output_if();
  logic c;
  modport port(output c);
endinterface: one_bit_output_if
