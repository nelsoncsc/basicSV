module hello();
  initial begin
    $display("hello from SV");
  end
endmodule
